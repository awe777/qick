module fixed_gauss(
	gauss_output,
);
output	[255:0]	gauss_output;
assign gauss_output = 256'h1337C0D3_DEADBEEF_CAFEBABE_0B00B135_4B1D4B1D_DEADC0DE_D0D0CACA_F0CACC1A;
endmodule